library IEEE;
use IEEE.std_logic_1164.ALL;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity symbol_rom is 
	port (	
		ADDRESS : in std_logic_vector(3 downto 0);
		COLUMN, ROW : in std_logic_vector(2 downto 0);
		DATA : out std_logic
	);
end symbol_rom;

architecture Behavioral of symbol_rom is
	type rom_array is array (0 to 15) of std_logic_vector(63 downto 0); 
	constant rom : rom_array := (
		"0000000000000000000000000000000000000000000000000000000000000000", -- prazdne policko?
		"0000000000010000000100000001000000010100000110000001000000000000", -- 1
		"0011110000000010000000100011110001000000010000000011110000000000", -- 2
		"0011110001000000010000000011100001000000010000000011110000000000", -- 3
		"0010000000100000001000000011111000100010001000100010001000000000", -- 4
		"0001111000100000001000000001110000000010000000100011110000000000", -- 5
		"0011110001000010010000100011110000000010000000100011110000000000", -- 6
		"0000010000000100000010000001000000100000001000000011111000000000", -- 7
		"0011110001000010010000100011110001000010010000100011110000000000", -- 8
		"0010000000100000001000000001110000100010001000100001110000000000", -- 9
		"0000000000110010010010100100101001001010010010100011001000000000", -- 10
		"0000000000100100001001000010010000100100001001000010010000000000", -- 11
		"0000000001110100000101000010010001000100010101000010010000000000", -- 12
		"0000000001110100010001000010010001000100010101000010000000000000", -- 13
		"0000000001000100010001000110010001010100010101000000000000000000", -- 14
		"0011100001000010010000100011001000001010000010100111001000000000"  -- 15
	);

begin
	result: process (ADDRESS, ROW, COLUMN) is
	begin
		data <= rom(conv_integer(ADDRESS))(conv_integer(ROW & COLUMN));
	end process result;
	
end Behavioral;

